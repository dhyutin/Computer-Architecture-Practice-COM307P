module testbench;
	reg s1, s2;
	reg [10:0] e1, e2;
	reg [51:0] m1, m2;
    
	wire [51:0] m;
	wire [10:0] e;
	wire s;
	
	dpfpm mult (s1, e1, m1, s2, e2, m2, s, m, e);

	initial begin
	    $dumpfile ("mult.vcd");
		$dumpvars (0,mult);
		s1 = 1'b0; e1 = 11'b10000000001; m1 = 52'b1100011001100110011001100110011001100110011001100110; 
		s2 = 1'b1; e2 = 11'b10000000010; m2 = 52'b0000011001100110011001100110011001100110011001100110; #10;

		s1 = 1'b1; e1 = 11'b10000000001; m1 = 52'b1100011001100110011001100110011001100110011001100110; 
		s2 = 1'b0; e2 = 11'b10000000010; m2 = 52'b0000011001100110011001100110011001100110011001100110; #10;
		
		s1 = 1'b0; e1 = 11'b10000000001; m1 = 52'b1100011001100110001101100010011001100110011001100110; 
		s2 = 1'b0; e2 = 11'b10000010010; m2 = 52'b0000011011110110001001100110011001100110011001100110; #10;
	end
	
	initial begin
		$monitor("\n s1 = %b, e1 = %b, m1 = %b, \n s2 = %b, e2 = %b, m2 = %b, \n s = %b, e = %b, m = %b,", s1, e1, m1, s2, e2, m2, s, e, m);  //$monitor is used to display the way form when the values change.
	end
endmodule